(** A simple module type for modules parameterized by a single
   type. *)
Module Type Sig.
Parameter A : Type.
End Sig.
